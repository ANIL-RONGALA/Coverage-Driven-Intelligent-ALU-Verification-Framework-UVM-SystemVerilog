//class 

class my_monitor extends uvm_monitor;
  `uvm_component_utils(my_monitor)
  
 
  virtual dut_if.MONITORPORT dut_vif_m;
  
  uvm_analysis_port#(my_transaction) monitor_ap;
  
  logic [31:0] in1_loc, in2_loc;
	op_e op_loc;

 
  //constructor
  function new(string name, uvm_component parent); 
    super.new(name, parent); 
    endfunction
      
    function void build_phase(uvm_phase phase); 
      //get interface reference from config database
        if(!uvm_config_db#(virtual dut_if.MONITORPORT)::get(this,"","dut_vif_m", dut_vif_m))  	
          begin
          `uvm_error("","uvm_config_db::get failed")
        end
      
      monitor_ap = new("monior_ap", this);
      
      endfunction
  
      
      // run phase 
      
      task run_phase(uvm_phase phase);
        my_transaction req;
      //check reset
         @(posedge dut_vif_m.clock);
        while(dut_vif_m.reset == 1)
          begin
            @(posedge dut_vif_m.clock);
       		 
          end
          @(posedge dut_vif_m.clock);
          @(posedge dut_vif_m.clock);
        @(posedge dut_vif_m.clock);
        in1_loc = dut_vif_m.in1;
        in2_loc = dut_vif_m.in2;
        op_loc = op_e'(dut_vif_m.cmd);
     
        forever begin
          
          @(posedge dut_vif_m.clock);
          req = my_transaction::type_id::create("req");
          
 		  req.in1 = in1_loc;
          req.in2 = in2_loc;
          req.op = op_loc;
          req.result = dut_vif_m.result;
          
          `uvm_info("MONITOR", $sformatf("Transaction generated by monitor - in1: %b, in2: %b, op: %h, result: = %b", req.in1, req.in2, req.op, req.result), UVM_LOW)
          
          monitor_ap.write(req);
          
          in1_loc = dut_vif_m.in1;
		  in2_loc = dut_vif_m.in2;
          op_loc = op_e'(dut_vif_m.cmd);
     
          
        
        end
          
      endtask

  
  endclass : my_monitor